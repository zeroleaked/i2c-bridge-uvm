`ifndef I2C_COMMON_PKG
`define I2C_COMMON_PKG

package i2c_common_pkg;
 
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	/////////////////////////////////////////////////////////
	// `include "i2c_interface.sv"

endpackage

`endif



