package i2c_master_wbs_8_pkg;
    import uvm_pkg::*;

	import i2c_common_pkg::*;

    // `include "sequence.svh"
    // `include "driver.svh"
    // `include "monitor.svh"
    // `include "agent.svh"
    // `include "scoreboard.svh"
    // `include "environment.svh"
    `include "test.svh"
endpackage