class write_read_seq extends uvm_sequence #(axil_seq_item);
    `uvm_object_utils(write_read_seq)
    
    function new(string name = "write_read_seq");
        super.new(name);
    endfunction

    task body();
        axil_seq_item req;
        bit [6:0] slave_addr = 7'h50;
        bit [7:0] reg_addr = 8'h0;
        bit [7:0] data_to_write = 8'hA5;
		
		memory_slave_seq mem_slave = memory_slave_seq::type_id::create("req");
		api_single_rw_seq api_rw = api_single_rw_seq::type_id::create("req");

		int timeout_count = 0;

        `uvm_info("SEQ", "Starting I2C write/read sequence", UVM_LOW)
        mem_slave.configure(m_sequencer, slave_addr);
		api_rw.configure(m_sequencer);
		
		mem_slave.register_write(reg_addr, data_to_write); // WRITE TO I2C SLAVE
        
        do begin
			api_rw.read_register_status();
            `uvm_info("SEQ", $sformatf("Status register: %h", api_rw.rsp.data), UVM_LOW)
        end while (api_rw.rsp.data[0]); // Wait until not busy
        
        #5000;
        
		// READ TO I2C SLAVE
		mem_slave.register_read(reg_addr);
        do begin
        	#100;
			timeout_count++;
			if (timeout_count > 10) begin
        		`uvm_error("SEQ", "Timeout waiting for a read")
				break;
			end
        end while (mem_slave.data[9:8] | DATA_VALID);
        
		`uvm_info("SEQ", $sformatf("Data register after read: %h", mem_slave.data), UVM_LOW)
    endtask
endclass