`ifndef I2C_AGENT_PKG
`define I2C_AGENT_PKG

package i2c_agent_pkg;
 
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	/////////////////////////////////////////////////////////

endpackage

`endif



